<!DOCTYPE html2
<head>
<title>Shasta System Management APIs</title>
<body>

  <h1>Shasta System Management Services</h1>

  <a href="l1/index.html">HaaS</a>
  <a href="l1/index.html">IaaS</a>
  <a href="l1/index.html">PaaS</a>


    <h2>Intro</h2>
    Intro
</body>
</html>


